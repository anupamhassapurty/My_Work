package mul_pkg;

	`include "transaction.sv"
	`include "sequence.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "agent.sv"
	`include "env.sv"
	`include "test.sv"

endpackage
