module tb;
    
	abp_if vif();
 
	apb_ram dut (vif.presetn, vif.pclk, vif.psel, vif.penable, vif.pwrite, vif.paddr, vif.pwdata, vif.prdata, vif.pready,vif.pslverr);
   
    initial begin
		vif.pclk <= 0;
    end
    
    always #10 vif.pclk <= ~vif.pclk;
    
    environment env;
     
    initial begin
		env = new(vif);
		env.gen.count = 30;
		env.run();
    end

    initial begin
      $dumpfile("dump.vcd");
      $dumpvars;
    end
   
endmodule
