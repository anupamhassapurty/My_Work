package add_pkg;

	`include "transaction.sv"
	`include "sequence1.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "agent.sv"
	`include "env.sv"
	`include "test.sv"

endpackage
