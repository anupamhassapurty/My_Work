interface add_if();
  logic clk;
  logic [3:0]a,b; 
  logic [3:0]sum;
  logic carry;
endinterface
