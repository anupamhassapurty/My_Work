interface mul_if;
	
	logic clk;	
	logic [7:0]m;
	logic [7:0]n;
	logic [15:0]mul;

endinterface
